module main

import json
import os

struct Patch {
  offset u64
  cleanbytes []u8
  patchbytes []u8
}
struct PatchScript{
 name string
 comment string
 patches []Patch
}

/*
commands
status patch_file infile
patch patch_file infile
clean patch_file infile
generate cleanfile patchfile
*/
	
       
fn main() {
  if os.args.len < 4 {
    println("Usage:\n ./PSOpatch status|patch|clean patch_file.json in_file.iso")
    return
  }
  match os.args[1] {
    'status' {
      patch_file := os.read_file(os.args[2])!
      test_file := os.open(os.args[3])!
      patch_script := json.decode(PatchScript, patch_file)!
      for patch in patch_script.patches {
	test_bytes := test_file.read_bytes_at(patch.patchbytes.len, patch.offset)
	  match test_bytes {
	    patch.cleanbytes {println("CLEAN")}
	    patch.patchbytes {println("PATCHED")}
	    else {println("MISMATCH")}
	  }
	}
    }
    'patch' {
      patch_file := os.read_file(os.args[2])!
      mut clean_file := os.open_file(os.args[3], 'r+')!
      patch_script := json.decode(PatchScript, patch_file)!
      for patch in patch_script.patches {
        clean_file.write_to(patch.offset, patch.patchbytes)!
      }
      clean_file.close()
    }
    'clean' {
      patch_file := os.read_file(os.args[2])!
      mut in_file := os.open_file(os.args[3], 'r+')!
      patch_script := json.decode(PatchScript, patch_file)!
      for patch in patch_script.patches {
        in_file.write_to(patch.offset, patch.cleanbytes)!
      }
      in_file.close()
    }
    'generate' {
      clean_file := os.open(os.args[2])!
      patch_file := os.open(os.args[3])!
      mut patches := []Patch{}
      mut offset := u64(0)
      mut in_patch := false
      mut patch_offset := u64(0)
      mut patch_clean := []u8{}
      mut patch_patch := []u8{}
      for clean_file.eof() == false && patch_file.eof() == false{      
        a := clean_file.read_bytes_at(1, offset)
        b := patch_file.read_bytes_at(1, offset)
        if a != b {
          if in_patch == false {
             in_patch = true
             patch_offset = offset
          }
          patch_clean << a
          patch_patch << b
        } else if in_patch {
          patches << Patch{patch_offset, patch_clean, patch_patch}
          in_patch = false
          patch_offset = 0
          patch_clean = []u8{}
          patch_patch = []u8{}
        }
        offset = offset + 1
      }
      patch_script := PatchScript{"Patch ${os.args[2]} to ${os.args[3]}", "Generated by PSOpatch", patches}
      println(json.encode_pretty(patch_script))
    }
    else {println("Unknown command!")}
  }

}
